* Circuito Modulador PWM por Doble Flanco para Audio

* Definici�n de componentes
.include LM741.MOD           ; Modelo de amplificador operacional LM741
.include LM393.MOD           ; Modelo de comparador LM393
.subckt TRIANG V+ V- OUT    ; Subcircuito para generador de onda triangular
R1 V+ 0 1k                   ; Resistencia de 1kO
R2 OUT V- 1k                 ; Resistencia de 1kO
C1 OUT 0 10u                 ; Capacitor de 10�F
.ends TRIANG

* Configuraci�n de componentes
Vmic IN 0 AC 1V SIN(0V 1V 1KHZ)     ; Fuente de audio (micr�fono simulado)
XOPAMP IN 0 OUT LM741              ; Amplificador operacional LM741
XTRI OUT 0 TRIANG                  ; Generador de onda triangular
XCOMP OUT 0 LM393                  ; Comparador LM393
RBNC OUT 0 50                      ; Carga resistiva para BNC

* An�lisis de transitorio
.TRAN 0.1MS 10MS                   ; An�lisis de transitorio de 0.1ms a 10ms

* Medici�n de variables
.PROBE
.END
