.TITLE Double-Edge PWM Modulator for Audio

* Define global simulation parameters
.OPTIONS TRAN 1uM 100m

* Define component models
.MODEL TIP41 NPN (BF=100)
.MODEL TIP31 PNP (BF=100)

* Define component values
R1 10k
R2 10k
R3 1k
R4 1k
R5 10k
C1 10u
C2 10u
C3 10u
C4 10u

* Define voltage sources
V1 5 0 DC 5V
V2 0 {AC 1V 1kHz} 

* Define 555 timer circuit
X1 1 2 3 4 5 6 7 8 555timer (VCC=V1 RST=0 TRIG=0)

* Define LM339 comparator circuit
X2 10 11 12 13 14 LM339 (VCC=V1 REF=V5 OUT=PWM)

* Define LM741 amplifier circuit
X3 15 16 17 18 19 LM741 (VCC=V1 VEE=0 IN=PWM OUT=AMP_PWM)

* Define TIP41 transistor circuit
Q1 20 21 22 TIP41 (VCC=V1 COLL=SPK BASE=AMP_PWM)

* Define speaker symbol
SPK 22 0 8

* Define BC547 transistor circuit
Q2 23 24 25 BC547 (VCC=V1 COLL=VCC BASE=V5)

* Define BC548 transistor circuit
Q3 26 27 28 BC548 (VCC=V1 COLL=VCC BASE=V2)

* Define potentiometer circuit
R6 29 30 10k
R7 30 0 10k

* Define voltage reference for LM339 comparator
V5 30 0 DC {LIN 0 5V 30k}

* Simulation output
.PROBE
.ENDP

.AC DEC 1 10k 100k
.END