.TITLE Double-Edge PWM Modulator for Audio

* Define component models
.MODEL TIP41 NPN (BF=100)
.MODEL TIP31 PNP (BF=100)

* Define component values
R1 10k
R2 10k
R3 1k
R4 1k
R5 10k
C1 10u
C2 10u
C3 10u
C4 10u

* Define voltage sources
V1 1 0 DC 5V
V2 2 0 SIN(0 1 1k)

* Define 555 timer circuit (replace with specific connections)
X1 1 2 3 4 5 6 7 8 555timer (VCC=V1 RST=0 TRIG=0)

* Define LM339 comparator circuit (replace with specific connections)
X2 9 10 11 12 13 LM339 (VCC=V1 REF=V5 OUT=PWM)

* Define LM741 amplifier circuit (replace with specific connections)
X3 14 15 16 17 18 LM741 (VCC=V1 VEE=0 IN=PWM OUT=AMP_PWM)

* Define TIP41 transistor circuit (replace with specific connections)
Q1 19 20 21 TIP41 (VCC=V1 COLL=SPK BASE=AMP_PWM)

* Define speaker symbol
SPK 20 0 8

* Define BC547 transistor circuit (replace with specific connections)
Q2 22 23 24 BC547 (VCC=V1 COLL=VCC BASE=V5)

* Define BC548 transistor circuit (replace with specific connections)
Q3 25 26 27 BC548 (VCC=V1 COLL=VCC BASE=V2)

* Define potentiometer circuit (replace with specific connections)
R6 28 29 10k
R7 29 0 10k

* Define voltage reference for LM339 comparator
V5 29 0 DC {LIN 0 5V 30k}

* Simulation output
.PROBE
.END

.AC DEC 1 10k 100k
.END