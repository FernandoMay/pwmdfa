* Double-Edge PWM Modulator for Audio

* Include Libraries
.include LM741.LIB
.include LM393.LIB
*.include 555.LIB
.MODEL 555 VCCS(RON=1G RS=1G)

* Micr�fono y Amplificador
Vmic IN 0 AC 1V SIN(0 1V 1kHz)
R1 IN 0 10k
C1 IN+ IN 10u
XOPAMP IN+ 0 OUT LM741
R4 OUT 0 10k

* Generador de Onda Triangular (555)
Vcc Vcc 0 DC 12V
X555 Vcc 0 0 TRIANG 555
R2 TRIANG Vcc 10k
R3 Vcc 0 4k7
C2 TRIANG 0 0.1u

* Comparador
XCOMP OUT+ TRIANG PWM LM393
R5 PWM 0 10k

* Amplificaci�n de la Se�al PWM
XAMP PWM 0 AMPOUT LM741
Q1 AMPOUT OUT1 Vcc TIP41
R6 OUT1 0 1k
RL OUT1 OUT2 8

* Salida
*BNC OUT2 0
*SPK OUT2 0

* Analysis
.TRAN 0.1ms 10ms
.PROBE
.END
