* PWM Modulation Circuit
* Generaci�n de Onda Triangular
*VCC 1 0 DC 12
*VEE 2 0 DC -12
R1 3 1 10k
C1 3 0 1uF
R2 3 4 10k
R3 4 2 10k
R4 4 0 10k
XU1 3 5 2 OPAMP
XU2 5 6 2 OPAMP
VTRI 6 0 SIN(0 1 1000)

* Comparadores
XU3 7 8 9 COMP
XU4 10 8 9 COMP
VAudio 8 0 SIN(0 1 100)
R5 7 0 10k
R6 10 0 10k

* Filtro Pasa-Bajos
R7 9 11 10k
C2 11 0 0.1uF

* Definici�n de Subcircuitos
.subckt OPAMP 1 2 3
* Pines: 1 = entrada positiva, 2 = entrada negativa, 3 = salida
E1 3 0 POLY(2) (1,2) (3,2) 1MEG
R1 3 0 10Meg
C1 3 0 1u
Rser 3 0 10
.ends OPAMP

.subckt COMP 1 2 3
* Pines: 1 = entrada positiva, 2 = entrada negativa, 3 = salida
E2 3 0 POLY(2) (1,2) (3,2) 1MEG
R2 3 0 10Meg
D1 3 0 D
.model D D
Rser 3 0 10
.ends COMP

* Fuentes de alimentaci�n
V1 1 0 DC 12
V2 2 0 DC -12

* Controles de simulaci�n
.tran 0.01ms 10ms
.end
